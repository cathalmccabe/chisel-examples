module Alu( // @[:@3.2]
  input  [1:0] io_fn, // @[:@6.4]
  input  [3:0] io_a, // @[:@6.4]
  input  [3:0] io_b, // @[:@6.4]
  output [3:0] io_result // @[:@6.4]
);
  wire  _T_16; // @[Conditional.scala 37:30:@10.4]
  wire [4:0] _T_17; // @[Alu.scala 37:27:@12.6]
  wire [3:0] _T_18; // @[Alu.scala 37:27:@13.6]
  wire  _T_20; // @[Conditional.scala 37:30:@17.6]
  wire [4:0] _T_21; // @[Alu.scala 38:27:@19.8]
  wire [4:0] _T_22; // @[Alu.scala 38:27:@20.8]
  wire [3:0] _T_23; // @[Alu.scala 38:27:@21.8]
  wire  _T_25; // @[Conditional.scala 37:30:@25.8]
  wire [3:0] _T_26; // @[Alu.scala 39:27:@27.10]
  wire  _T_28; // @[Conditional.scala 37:30:@31.10]
  wire [3:0] _T_29; // @[Alu.scala 40:27:@33.12]
  wire [3:0] _GEN_0; // @[Conditional.scala 39:67:@32.10]
  wire [3:0] _GEN_1; // @[Conditional.scala 39:67:@26.8]
  wire [3:0] _GEN_2; // @[Conditional.scala 39:67:@18.6]
  assign _T_16 = 2'h0 == io_fn; // @[Conditional.scala 37:30:@10.4]
  assign _T_17 = io_a + io_b; // @[Alu.scala 37:27:@12.6]
  assign _T_18 = _T_17[3:0]; // @[Alu.scala 37:27:@13.6]
  assign _T_20 = 2'h1 == io_fn; // @[Conditional.scala 37:30:@17.6]
  assign _T_21 = io_a - io_b; // @[Alu.scala 38:27:@19.8]
  assign _T_22 = $unsigned(_T_21); // @[Alu.scala 38:27:@20.8]
  assign _T_23 = _T_22[3:0]; // @[Alu.scala 38:27:@21.8]
  assign _T_25 = 2'h2 == io_fn; // @[Conditional.scala 37:30:@25.8]
  assign _T_26 = io_a | io_b; // @[Alu.scala 39:27:@27.10]
  assign _T_28 = 2'h3 == io_fn; // @[Conditional.scala 37:30:@31.10]
  assign _T_29 = io_a & io_b; // @[Alu.scala 40:27:@33.12]
  assign _GEN_0 = _T_28 ? _T_29 : 4'h0; // @[Conditional.scala 39:67:@32.10]
  assign _GEN_1 = _T_25 ? _T_26 : _GEN_0; // @[Conditional.scala 39:67:@26.8]
  assign _GEN_2 = _T_20 ? _T_23 : _GEN_1; // @[Conditional.scala 39:67:@18.6]
  assign io_result = _T_16 ? _T_18 : _GEN_2; // @[Alu.scala 44:13:@36.4]
endmodule
module AluTop( // @[:@38.2]
  input        clock, // @[:@39.4]
  input        reset, // @[:@40.4]
  input  [9:0] io_sw, // @[:@41.4]
  output [9:0] io_led // @[:@41.4]
);
  wire [1:0] alu_io_fn; // @[Alu.scala 57:19:@43.4]
  wire [3:0] alu_io_a; // @[Alu.scala 57:19:@43.4]
  wire [3:0] alu_io_b; // @[Alu.scala 57:19:@43.4]
  wire [3:0] alu_io_result; // @[Alu.scala 57:19:@43.4]
  Alu alu ( // @[Alu.scala 57:19:@43.4]
    .io_fn(alu_io_fn),
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_result(alu_io_result)
  );
  assign io_led = {{6'd0}, alu_io_result}; // @[Alu.scala 65:10:@52.4]
  assign alu_io_fn = io_sw[1:0]; // @[Alu.scala 60:13:@47.4]
  assign alu_io_a = io_sw[5:2]; // @[Alu.scala 61:12:@49.4]
  assign alu_io_b = io_sw[9:6]; // @[Alu.scala 62:12:@51.4]
endmodule
